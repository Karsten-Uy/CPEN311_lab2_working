// TODO: see if this needs to be in a seperate file or could just be
// in the package

interface phases;

    logic reset_phase;
    logic run_phase;
    logic report_phase;
    
endinterface // phases

