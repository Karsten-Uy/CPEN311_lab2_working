interface phases;

    logic reset_phase;
    logic run_phase;
    logic report_phase;
    
endinterface // phases

