interface top_if ;

    logic           CLOCK_50;
    logic   [3:0]   KEY;
    logic   [9:0]   LEDR;
    logic   [6:0]   HEX5;
    logic   [6:0]   HEX4;
    logic   [6:0]   HEX3;
    logic   [6:0]   HEX2;
    logic   [6:0]   HEX1;
    logic   [6:0]   HEX0;
    
endinterface //datapath_if

